------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
------------

entity DrinksFSMTB is
			
end DrinksFSMTB;
-------------

architecture Silva of DrinksFSM is
	type state_type is(S0, S1, S2, S3, S4, S5, S6, S7);
	Signal s_pstate, state_next : state_type;
begin
		
end Silva;
---------