---------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
---------------

entity ALU4 is
			port(a, b : in std_logic_vector(3 downto 0);
				 op 	 : in std_logic_vector(2 downto 0);
				 r, m  : out std_logic_vector(3 downto 0));
end ALU4;
--------------

architecture Behavioral of ALU4 is

	signal s_a, s_b, s_r : signed(3 downto 0);
	signal s_m           : signed(7 downto 0);
	
begin
				 s_a <= signed(a);
				 s_b <= signed(b);
				 s_m <= s_a * s_b; 
				 
				
				 s_r <= s_a + s_b         when (op = "000") else
						  s_a - s_b         when (op = "001") else
						  s_m(3 downto 0)   when (op = "010") else
						  s_a / s_b   		  when (op = "011") else
						  s_a rem s_b       when (op = "100") else
						  s_a and s_b       when (op = "101") else
						  s_a or s_b  		  when (op = "110") else
						  s_a xor s_b       when (op = "111");
				 r <= std_logic_vector(s_r);
				 m <= std_logic_vector(s_m(7 downto 4)) when (op = "010") else
				 (others => '0');
end Behavioral;
--------------