------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
------------

entity cntUp is
				port(clk 	: in std_logic;
					  reset  : in std_logic;
					  enable : in std_logic;
					  cntval : out std_logic_vector(29 downto 0));
end cntup;
---------

architecture behavioral of cntup is 
	signal s_cntup : unsigned(29 downto 0);
	
begin 
		
		process(clk)
			begin
				 if(rising_edge(clk)) then 
					if(reset = '1') then 
						s_cntup <= (others => '0');
						
					 elsif(enable = '1') then 
						s_cntup <= s_cntup + 1;
						
					end if;
				 end if;
			end process;
	cntval <= std_logic_vector(s_cntup);
	
end behavioral;
			